Differentiator
*Including the predefined op-amp subcircuit file
.include uA741.txt

C1 1 2 0.01u
VCC 4 gnd dc 15
VEE 5 gnd dc -15
x1 gnd 2 4 5 3 uA741
R1 2 3 10k
C2 2 3 0.001u
Vi 1 gnd pulse(-2 2 0 0.2m 0.2m 1n 0.4m)

.tran 0.00005m 3m
.control
run

plot v(1) v(3)

.endc
.end
