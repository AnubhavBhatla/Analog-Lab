RC Bandpass Filter

*Connections as mentioned in the subcircuit file
R1 1 2 10k
C1 2 3 0.1u
R2 3 0 10k
C2 3 0 0.1u

*Giving an input
Vin 1 0 dc 0 ac 1

.ac dec 1000 1 1Meg
.control
run

plot vdb(3)
print vdb(3)
.endc
.end
