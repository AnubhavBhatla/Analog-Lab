Inverting Schmitt Trigger
*Including the predefined subcircuit files
.include zener_1N4732A.txt
.include ua741.txt
.include Diode_1N914.txt

R1 5 2 13.3k
R2 6 3 13.3k
VCC 5 0 dc 15
VEE 6 0 dc -15
x1 out in 5 6 out ua741
D1 2 1 1N914
D2 2 out 1N914
D3 1 3 1N914
D4 out 3 1N914
x2 out 4 DI_1N4732A
x3 0 4 DI_1N4732A
Vin in 0 sin(0 6 1k 0 0)

.tran 0.01m 5m

.control
run

plot v(out) v(in)

.endc
.end
