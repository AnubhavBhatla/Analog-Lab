Inverting Schmitt Trigger
*Including the predefined subcircuit files
.include zener_1N4732A.txt
.include ua741.txt
.include Diode_1N914.txt

R1 5 2 13.3k
R2 6 3 13.3k
VCC 5 0 dc 15
VEE 6 0 dc -15
x1 out in 5 6 out ua741
D1 2 1 1N914
D2 2 out 1N914
D3 1 3 1N914
D4 out 3 1N914
x2 out 4 DI_1N4732A
x3 0 4 DI_1N4732A
Vin in 0 dc 0

.control

dc Vin 10 -10 -0.1

*dc Vin -10 10 0.1

plot v(out) 

.endc
.end
