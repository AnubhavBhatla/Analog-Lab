Circuit - 3a
*Including the predefined op-amp subcircuit file
.include zener_B.txt
.include uA741.txt

R1 1 2 8.2k
R2 2 3 15k
R3 4 3 1k
VCC 5 0 dc 15
VEE 6 0 dc -15
x1 2 0 5 6 4 uA741
x2 3 7 DI_1N4734A
x3 0 7 DI_1N4734A
Vin 1 0 dc 0

.dc Vin -5 5 0.01
.control
run

plot v(3)

.endc
.end
