RC Differentiator

*Connections as mentioned in the subcircuit file
C 1 2 0.1u
R 2 0 10k

*Giving an input
Vin 1 0 pulse(0 5 0 0 0 10m 20m)

.tran 0.02m 60m
.control
run

plot v(1) v(2)
print v(1) v(2)
.endc
.end
