Circuit - 2
*Including the predefined op-amp subcircuit file
.include uA741.txt

Rx1 1 2 10k
Rx2 2 4 10k
R 1 3 1k
C 3 0 1n
VCC 5 0 dc 15
VEE 6 0 dc -15
x1 3 2 5 6 4 uA741
Vi 1 0 dc 0 ac 0.5

.ac dec 100 1 1Meg
.control
run

plot {20*log(v(4)/v(1))}
plot {57.29*vp(4)}

.endc
.end
