Bridge Rectifier

*Model file for the Diode
.MODEL 1N4007 D (IS=76.9p RS=42.0m BV=1k IBV=1
+ CJO=26.5p  M=0.333 N=1.45 TT=4.32u)

d1 dummy1 2 1N4007
d2 0 1 1N4007
d3 dummy3 2 1N4007
d4 0 3 1N4007
Rl 2 0 1k
Vd1 1 dummy1 dc 0
Vd2 3 dummy3 dc 0
Vin 1 3 sin(0 21.21 50 0 0)

.tran 0.1m 100m
.control
run

plot v(2)
plot i(Vd1) i(Vd2)

.endc
.endA
