RLC Bandpass Filter

*Connections as mentioned in the subcircuit file
L 1 2 10m
C 2 3 0.1u
R 3 0 1k

*Giving an input
Vin 1 0 dc 0 ac 1

.ac dec 100 1 1Meg
.control
run

plot vdb(3)
print vdb(3)
.endc
.end
