Wheat-Stone Bridge
*Including the predefined op-amp subcircuit file
.include lm324.txt

Ra 1 0 300
Rc 2 1 300
Rb 2 3 300
Rx 3 0 300
R1 3 4 2.5k
R2 4 0 100k
R3 5 6 100k
R4 6 1 2.5k
VCC 7 0 dc 15
VEE 8 0 dc -15
x1 4 6 7 8 5 LM324
V1 2 0 dc 5

.dc Rx 300 310 5
.control
run

plot v(1,3)
plot v(5)

.endc
.end
