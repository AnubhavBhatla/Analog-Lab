Wheat-Stone Bridge with Thermistor
*Including the predefined subcircuit files
.include lm324.txt
.include Thermistor.txt

Ra 1 0 300
Rc 2 1 300
Rb 2 3 300
x2 3 0 9 thermistor Ro=300 alpha=-3548  
R1 3 4 2k
R2 4 0 10k
R3 5 6 10k
R4 6 1 2k
VCC 7 0 dc 15
VEE 8 0 dc -15
x1 4 6 7 8 5 LM324
V1 2 0 dc 5
Vtemp 9 0 dc 0

.dc Vtemp 20 30 0.1
.control
run

plot v(1,3)
plot v(5)

.endc
.end
