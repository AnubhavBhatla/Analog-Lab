Unregulated Supply

*Model file for the Diode
.MODEL 1N4007 D (IS=76.9p RS=42.0m BV=1k IBV=1
+ CJO=26.5p  M=0.333 N=1.45 TT=4.32u)

.param cap=100u

d1 1 2 1N4007
d2 0 1 1N4007
d3 3 2 1N4007
d4 0 3 1N4007
Rl 2 0 500
C1 2 0 cap
Vin 1 3 sin(0 21.21 50 0 0)

.control

alter C1=100u
tran 0.01m 100m

alter C1=470u
tran 0.01m 100m

alter C1=1000u
tran 0.01m 100m

plot tran1.v(2) tran2.v(2) tran3.v(2)
.endc
.end
