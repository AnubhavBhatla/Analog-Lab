Circuit 2-c
*Including the predefined subcircuit files
.include lm324.txt

RG in 1 8.2k
RF 1 out 120k
R1 2 0 8.2k
R2 ref 2 120k
Vref ref 0 10.4
VCC 3 0 dc 5
VEE 4 0 dc 0
x1 2 1 3 4 out lm324
Vin in 0 dc 0

.dc Vin 0 2 0.01
.control
run

plot v(out) vs v(in)

.endc
.end
