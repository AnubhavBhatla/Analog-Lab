Full-Wave Precision Rectifier
*Including the predefined op-amp subcircuit file
.include HWPR_B_S.txt
.include uA741.txt

x1 1 2 HWPR
R1 1 3 10k
R2 2 3 5k
R3 3 4 10k
Rl 4 0 1k
VCC 5 0 dc 15
VEE 6 0 dc -15
x2 0 3 5 6 4 uA741
Vi 1 0 sin(0 5 1k 0 0)

.tran 0.0001m 4m
.control
run

print v(4) v(1)

.endc
.end
