Photodiode
*Including the predefined subcircuit files
.include lm324.txt

I1 1 0 0
CJ 1 0 11p
x1 2 1 4 5 out lm324
R1 1 out 1.4Meg
C1 1 out 3.3p
R2 2 4 13.7k
R3 2 0 280
C2 2 0 1u
Vref 2 0 dc 0.1
VCC 4 0 dc 5
VEE 5 0 dc 0

.dc I1 0 2.4u 0.1u
.control
run

plot v(out)

.endc
.end
