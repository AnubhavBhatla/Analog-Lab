Half-Wave Precision Rectifier - B
*Including the predefined op-amp subcircuit file
.include uA741.txt

R1 1 2 10k
R2 2 3 10k
Rl 3 0 1k
D1 4 2
D2 3 4
VCC 5 0 dc 15
VEE 6 0 dc -15
x1 0 2 5 6 4 uA741
Vi 1 0 sin(0 5 1k 0 0)

.tran 0.0001m 4m
.control
run

print v(1) v(3) v(4)

.endc
.end
